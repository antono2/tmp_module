module tmp_module

pub const v_modroot = @VMODROOT
