module tmp_module

pub const v_modroot = @VMODROOT

pub struct MyParentStruct{
pub mut:
  value int
}

