module another_module

pub const v_modroot = @VMODROOT
